

//preset the rx, because idle is high, and start bit is low